module Sample(